`timescale 1ns/1ps
`default_nettype none

module tb_uart_harness(
    inout wire rx
);
endmodule